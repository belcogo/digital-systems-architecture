module behav_and_gate (A, B, S);
    input A, B;
    output S;

    assign S = A & B;
endmodule